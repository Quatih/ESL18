-- QuadDec.vhd

-- Generated using ACDS version 13.0sp1 232 at 2018.05.18.14:15:25

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity QuadDec is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity QuadDec;

architecture rtl of QuadDec is
begin

end architecture rtl; -- of QuadDec
